library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY SSegment IS									
	PORT(					
        CLK      :  IN STD_LOGIC;   
				BCD_In   :  IN STD_LOGIC_VECTOR(3 DOWNTO 0);	
				Segment  : 	OUT STD_LOGIC_VECTOR(6 DOWNTO 0)			
		);																	
END SSegment;
--------------------------------------------------------------------
--                 Architecture of SSegment
--------------------------------------------------------------------

ARCHITECTURE Beh_SSegment OF SSegment IS			-- Counter = Entity Name
	signal SegmentInt  :  STD_LOGIC_VECTOR(6 DOWNTO 0)	;
BEGIN

   WITH BCD_In SELECT					-- Auswahl
	Segment  <= "1000000" WHEN x"0",
		      "1111001" WHEN x"1",		--	    0			 
		      "0100100" WHEN x"2",		--	   ---
		      "0110000" WHEN x"3",		--	 5| 6 |1
		      "0011001" WHEN x"4",		--	   ---
		      "0010010" WHEN x"5",		--	 4|   |2
		      "0000010" WHEN x"6",		--	   ---
		      "1111000" WHEN x"7",		--	    3
		      "0000000" WHEN x"8",
		      "0010000" WHEN x"9",
		      "1111111" WHEN OTHERS;   

END Beh_SSegment;
