-- A library clause declares a name as a library.  It 
-- does not create the library; it simply forward declares 
-- it. 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_signed.all;

-- Library Clause(s) (optional)
-- Use Clause(s) (optional)
entity Game_Main is

	port
	(
		-- Input ports
			xpos_game     					:	in  	integer range 0 to 1300;   						-- Pixel Pos x Bildbereich
			ypos_game     					:	in  	integer range 0 to 1033;    					-- Pixel Pos y Bildbereich
			BTN_LEFT								:	in	 	std_logic;
			BTN_RIGHT								:	in	 	std_logic;
			Reset										:	in		std_logic;
			videoOn_game  					:	in  	std_logic;               							-- 1 = Bildbereich
			vga_clk									:	in		std_logic;
			NewFrame_game						:	in		std_logic;	

		-- Inout ports


		-- Output ports
			Draw_Snake_Out							: out 	std_logic := 	'0';
			Draw_Apple_Out							:	out		std_logic	:=	'0');
end Game_Main;

architecture beh_Game_Main of Game_Main is

	-- Declarations (optional)
	-- Signal Declarations
	
	signal 			Draw_Apple_In							:	std_logic	:= '0';
	signal 			Draw_Snake_In							:	std_logic	:= '0';
	signal 			Add												:	std_logic	:= '0';
	signal			x_Apple_Game							:	integer range	0	to	2000 := 0;
	signal			y_Apple_Game							:	integer range	0	to	2000 := 0;
	signal			x_snake_Game							:	integer range	0	to	2000 := 0;
	signal			y_snake_Game							:	integer range	0	to	2000 := 0;

begin

	/*Snake_Drawing Instantiation*/
		
		Snake_Drawing	:	entity	work.snake_Drawing
			port map (
					xpos_snake     					=>	xpos_game,
					ypos_snake     					=>	ypos_game,
					BTN_LEFT								=>	BTN_LEFT,
					BTN_RIGHT								=>	BTN_RIGHT,
					videoOn_snake  					=>	videoOn_game,
					vga_clk									=>	vga_clk,
					NewFrame_snake					=>	NewFrame_game,
					Draw_Snake							=>	Draw_Snake_In,
					Reset										=>	Reset,
					x_pos_snake						=>	x_snake_Game,
					y_pos_snake						=>	y_snake_Game,
					add_snake								=>	add);
					
	/*Apple_Drawing Instantiation*/
		Apple_Drawing	: entity	work.Apple_Drawing
			port map(
					xpos_apple     					=>	xpos_game,
					ypos_apple     					=>	ypos_game,
					videoOn_apple  					=>	videoOn_game,
					vga_clk									=>	vga_clk,
					NewFrame_apple					=>	NewFrame_game,
					Draw_apple							=>	Draw_Apple_In,
					Reset										=>	Reset,
					x_Apple_OUT							=>	x_apple_Game,
					y_apple_Out							=>	y_apple_Game
			);
			
					
				Game_Main : process(all)
				
				begin
						
						if rising_edge(vga_clk)	then
							
							Draw_Apple_Out <= Draw_Apple_In;
							Draw_Snake_Out <=	Draw_Snake_In;
							
							if x_apple_Game = x_snake_Game and y_apple_Game = y_snake_Game	then
								Add <= '1';
							else
								Add <= '0';
							end if;
							
							
						end if;
						
				end process Game_Main;
	-- Process Statement (optional)

	-- Concurrent Procedure Call (optional)

	-- Concurrent Signal Assignment (optional)

	-- Conditional Signal Assignment (optional)

	-- Selected Signal Assignment (optional)

	-- Component Instantiation Statement (optional)

	-- Generate Statement (optional)

end beh_Game_Main;

